bind dma dma_checker_sva check1(busIf);
bind dma dma_checker_sva_reset check2(busIf);
