bind dma dma_checker_sva check1(busIf);
