bind dma dma_checker_sva_eop check3(busIf);
