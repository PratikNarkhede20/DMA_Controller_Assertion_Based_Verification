bind dma dma_checker_sva_reset check2(busIf);
