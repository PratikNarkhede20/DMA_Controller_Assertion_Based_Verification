bind dma dma_checker_sva_run check1(busIf);
