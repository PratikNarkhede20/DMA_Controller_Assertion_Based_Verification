module dma_checker_sva(busInterface busIf);


default clocking c0 @(posedge busIf.CLK); endclocking



endmodule
